`timescale 1us / 1ps
